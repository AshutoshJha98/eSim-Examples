* /home/ash98/Downloads/eSim-master/src/SubcircuitLibrary/Ideal_OpAmp/Ideal_OpAmp.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Tue Dec 31 11:36:29 2019

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
Q3  Net-_Q2-Pad1_ Net-_Q2-Pad1_ Net-_Q3-Pad3_ eSim_PNP		
Q5  Net-_C1-Pad2_ Net-_Q2-Pad1_ Net-_Q3-Pad3_ eSim_PNP		
Q2  Net-_Q2-Pad1_ /Inv Net-_Q2-Pad3_ eSim_NPN		
Q6  Net-_C1-Pad2_ /Non-Inv Net-_Q2-Pad3_ eSim_NPN		
Q4  Net-_Q2-Pad3_ Net-_Q1-Pad1_ Net-_Q1-Pad3_ eSim_NPN		
Q1  Net-_Q1-Pad1_ Net-_Q1-Pad1_ Net-_Q1-Pad3_ eSim_NPN		
R1  Net-_Q3-Pad3_ Net-_Q1-Pad1_ 9.8k		
R2  Net-_Q3-Pad3_ Net-_D1-Pad1_ 5.11k		
Q7  Net-_C1-Pad1_ Net-_C1-Pad2_ Net-_Q3-Pad3_ eSim_PNP		
D1  Net-_D1-Pad1_ Net-_D1-Pad2_ eSim_Diode		
C1  Net-_C1-Pad1_ Net-_C1-Pad2_ 400p		
R3  Net-_D1-Pad2_ Net-_Q1-Pad3_ 20		
Q8  Net-_C1-Pad1_ Net-_D1-Pad1_ Net-_Q1-Pad3_ eSim_NPN		
Q9  Net-_Q3-Pad3_ Net-_C1-Pad1_ /Out eSim_NPN		
Q10  /Out Net-_D1-Pad1_ Net-_Q1-Pad3_ eSim_NPN		
U1  /Inv /Non-Inv /Out Net-_Q3-Pad3_ Net-_Q1-Pad3_ PORT		

.end
