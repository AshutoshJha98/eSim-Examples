* /home/ash98/Downloads/eSim-master/src/SubcircuitLibrary/Ideal_OpAmp/Ideal_OpAmp.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Sat Dec 28 17:17:21 2019

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
Q4  Net-_C1-Pad2_ Net-_Q2-Pad1_ Net-_Q13-Pad1_ eSim_NPN		
Q1  GND /Inv Net-_Q1-Pad3_ eSim_PNP		
Q2  Net-_Q2-Pad1_ Net-_Q1-Pad3_ Net-_Q2-Pad3_ eSim_PNP		
Q6  GND /Non-Inv Net-_Q5-Pad2_ eSim_PNP		
Q5  Net-_C1-Pad2_ Net-_Q5-Pad2_ Net-_Q2-Pad3_ eSim_PNP		
Q3  Net-_Q13-Pad1_ Net-_Q2-Pad1_ Net-_Q2-Pad1_ eSim_NPN		
Q11  Net-_Q11-Pad1_ Net-_C1-Pad1_ Net-_Q11-Pad3_ eSim_NPN		
Q12  Net-_Q11-Pad1_ Net-_Q11-Pad3_ Net-_Q10-Pad2_ eSim_NPN		
Q13  Net-_Q13-Pad1_ Net-_C1-Pad1_ /Out eSim_PNP		
Q10  Net-_C1-Pad1_ Net-_Q10-Pad2_ /Out eSim_NPN		
Q8  Net-_Q8-Pad1_ Net-_Q7-Pad3_ Net-_Q8-Pad3_ eSim_NPN		
Q9  Net-_C1-Pad1_ Net-_Q8-Pad3_ Net-_Q13-Pad1_ eSim_NPN		
Q7  ? Net-_C1-Pad2_ Net-_Q7-Pad3_ eSim_PNP		
U1  /Inv /Non-Inv /Out Net-_Q11-Pad1_ Net-_Q13-Pad1_ PORT		
C1  Net-_C1-Pad1_ Net-_C1-Pad2_ 50p		
R2  Net-_Q10-Pad2_ /Out 30		
R1  Net-_Q8-Pad3_ Net-_Q13-Pad1_ 100k		
R3  Net-_Q11-Pad1_ Net-_Q2-Pad3_ 300k		
R4  Net-_Q11-Pad1_ Net-_Q8-Pad1_ 500k		
R5  Net-_Q11-Pad1_ Net-_C1-Pad1_ 50k		
R6  /Out Net-_Q13-Pad1_ 100k		

.end
