* /home/ash98/eSim-Workspace/Ina128/Ina128.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Sat Dec 28 10:10:49 2019

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
X1  Net-_R3-Pad1_ Net-_R1-Pad2_ GND Net-_X1-Pad4_ GND Out Net-_X1-Pad7_ Net-_R3-Pad2_ INA_128		
v1  In GND sine		
R1  In Net-_R1-Pad2_ 1k		
R3  Net-_R3-Pad1_ Net-_R3-Pad2_ 1k		
R4  Out GND 1k		
v3  Net-_X1-Pad7_ GND DC		
v2  GND Net-_X1-Pad4_ DC		
R2  Net-_R1-Pad2_ Out 10k		
U1  In plot_v1		
U2  Out plot_v1		

.end
