* /home/ash98/Downloads/LM_386N/LM_386N.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Fri Dec 27 13:26:08 2019

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
Q3  Net-_Q2-Pad1_ Net-_Q2-Pad1_ /Gnd eSim_NPN		
Q2  Net-_Q2-Pad1_ Net-_Q1-Pad3_ Net-_Q2-Pad3_ eSim_PNP		
R2  /Vcc Net-_R2-Pad2_ 15k		
R3  Net-_R2-Pad2_ Net-_Q2-Pad3_ 15k		
U1  Net-_Q5-Pad3_ Net-_Q1-Pad2_ Net-_Q6-Pad2_ /Gnd /Out /Vcc Net-_R2-Pad2_ Net-_R4-Pad1_ PORT		
R4  Net-_R4-Pad1_ Net-_Q2-Pad3_ 150		
R5  Net-_Q5-Pad3_ Net-_R4-Pad1_ 1.35k		
Q5  Net-_Q4-Pad1_ Net-_Q5-Pad2_ Net-_Q5-Pad3_ eSim_PNP		
R7  /Out Net-_Q5-Pad3_ 15k		
Q1  /Gnd Net-_Q1-Pad2_ Net-_Q1-Pad3_ eSim_PNP		
R1  Net-_Q1-Pad2_ /Gnd 50k		
Q4  Net-_Q4-Pad1_ Net-_Q2-Pad1_ /Gnd eSim_NPN		
Q6  /Gnd Net-_Q6-Pad2_ Net-_Q5-Pad2_ eSim_PNP		
R6  Net-_Q6-Pad2_ /Gnd 50k		
Q7  Net-_D2-Pad2_ Net-_Q4-Pad1_ /Gnd eSim_NPN		
D1  Net-_D1-Pad1_ Net-_D1-Pad2_ eSim_Diode		
D2  Net-_D1-Pad2_ Net-_D2-Pad2_ eSim_Diode		
Q9  /Vcc Net-_D1-Pad1_ /Out eSim_NPN		
Q10  /Out Net-_Q10-Pad2_ /Gnd eSim_NPN		
Q8  Net-_Q10-Pad2_ Net-_D2-Pad2_ /Out eSim_PNP		
R8  /Vcc Net-_D1-Pad1_ 10k		

.end
