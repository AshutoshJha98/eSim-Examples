* /home/ash98/Downloads/eSim-master/src/SubcircuitLibrary/MPY_634/MPY_634.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Tue Dec 31 16:55:23 2019

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U3  Net-_U1-Pad3_ Net-_U2-Pad3_ Net-_U3-Pad3_ mult		
U5  Net-_U3-Pad3_ Net-_U5-Pad2_ Net-_U5-Pad3_ divide		
U1  Net-_R3-Pad2_ Net-_U1-Pad2_ Net-_U1-Pad3_ summer		
U2  Net-_R4-Pad2_ Net-_U2-Pad2_ Net-_U2-Pad3_ summer		
U6  Net-_R6-Pad2_ Net-_U6-Pad2_ Net-_U6-Pad3_ summer		
U8  Net-_U1-Pad2_ Net-_R1-Pad1_ ? Net-_U5-Pad2_ ? Net-_U2-Pad2_ Net-_R2-Pad1_ Net-_U8-Pad8_ ? Net-_U6-Pad2_ Net-_R5-Pad1_ Net-_U4-Pad2_ ? /+Vs PORT		
U9  Net-_U6-Pad3_ Net-_U5-Pad3_ Net-_U4-Pad1_ summer		
X1  Net-_R1-Pad2_ GND Net-_R3-Pad2_ /+Vs Net-_U8-Pad8_ OpAmp_1		
X2  Net-_R2-Pad2_ GND Net-_R4-Pad2_ /+Vs Net-_U8-Pad8_ OpAmp_1		
X3  Net-_R5-Pad2_ GND Net-_R6-Pad2_ /+Vs Net-_U8-Pad8_ OpAmp_1		
R1  Net-_R1-Pad1_ Net-_R1-Pad2_ 1k		
R3  Net-_R1-Pad2_ Net-_R3-Pad2_ 1k		
R2  Net-_R2-Pad1_ Net-_R2-Pad2_ 1k		
R4  Net-_R2-Pad2_ Net-_R4-Pad2_ 1k		
R5  Net-_R5-Pad1_ Net-_R5-Pad2_ 1k		
R6  Net-_R5-Pad2_ Net-_R6-Pad2_ 1k		
U4  Net-_U4-Pad1_ Net-_U4-Pad2_ gain		

.end
