* /home/ash98/Downloads/eSim-master/src/SubcircuitLibrary/INA_128/INA_128.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Fri Dec 27 16:51:24 2019

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
X1  ? Net-_R1-Pad1_ /-Vin Net-_U1-Pad4_ ? Net-_R1-Pad2_ Net-_U1-Pad7_ ? lm_741		
X2  ? Net-_R2-Pad1_ /+Vin Net-_U1-Pad4_ ? Net-_R2-Pad2_ Net-_U1-Pad7_ ? lm_741		
X3  ? Net-_R3-Pad2_ Net-_R4-Pad2_ Net-_U1-Pad4_ ? Net-_R5-Pad2_ Net-_U1-Pad7_ ? lm_741		
R1  Net-_R1-Pad1_ Net-_R1-Pad2_ 25k		
R2  Net-_R2-Pad1_ Net-_R2-Pad2_ 25k		
R4  Net-_R2-Pad2_ Net-_R4-Pad2_ 40k		
R3  Net-_R1-Pad2_ Net-_R3-Pad2_ 40k		
R5  Net-_R3-Pad2_ Net-_R5-Pad2_ 40k		
R6  Net-_R4-Pad2_ /Ref 40k		
U1  Net-_R1-Pad1_ /-Vin /+Vin Net-_U1-Pad4_ /Ref Net-_R5-Pad2_ Net-_U1-Pad7_ Net-_R2-Pad1_ PORT		

.end
