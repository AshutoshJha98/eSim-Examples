* /home/ash98/eSim-Workspace/Therm2binary/Therm2binary.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Fri Jan  3 15:09:12 2020

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U2  Ref2 plot_v1		
U3  Ref3 plot_v1		
U1  Ref1 plot_v1		
X1  ? Net-_R5-Pad1_ Net-_R6-Pad1_ Net-_X1-Pad4_ ? Out1 Net-_X1-Pad7_ ? lm_741		
R5  Net-_R5-Pad1_ Ref1 1k		
X2  ? Net-_R7-Pad1_ Net-_R8-Pad1_ Net-_X1-Pad4_ ? Out2 Net-_X1-Pad7_ ? lm_741		
R7  Net-_R7-Pad1_ Ref2 1k		
X3  ? Net-_R9-Pad1_ Net-_R10-Pad1_ Net-_X1-Pad4_ ? Out3 Net-_X1-Pad7_ ? lm_741		
R9  Net-_R9-Pad1_ Ref3 1k		
R6  Net-_R6-Pad1_ V_In 1k		
R8  Net-_R8-Pad1_ V_In 1k		
R10  Net-_R10-Pad1_ V_In 1k		
R11  Net-_R11-Pad1_ Out1 1k		
R12  Net-_R12-Pad1_ Out2 1k		
R13  Net-_R13-Pad1_ Out3 1k		
v3  Net-_X1-Pad7_ GND 6		
U4  Out1 plot_v1		
U5  Out2 plot_v1		
U6  Out3 plot_v1		
v4  GND Net-_X1-Pad4_ 6		
U7  Net-_R11-Pad1_ Net-_R12-Pad1_ Net-_R13-Pad1_ Net-_U7-Pad4_ Net-_U7-Pad5_ Net-_U7-Pad6_ adc_bridge_3		
U9  Net-_U8-Pad4_ Net-_U8-Pad5_ Bin1 Bin2 dac_bridge_2		
R15  GND Bin1 1k		
R14  Bin2 GND 1k		
U11  Bin1 plot_v1		
U10  Bin2 plot_v1		
U12  V_In plot_v1		
v1  Net-_R1-Pad2_ GND 4		
R1  Ref1 Net-_R1-Pad2_ 1k		
R2  Ref2 Ref1 1k		
R3  Ref3 Ref2 1k		
R4  GND Ref3 1k		
v2  V_In GND DC		
U8  Net-_U7-Pad4_ Net-_U7-Pad5_ Net-_U7-Pad6_ Net-_U8-Pad4_ Net-_U8-Pad5_ therm2bin2bit		

.end
